    /*
     * Small Vector Floating Point RISC-V Core
     *
     * @copyright 2025 Paolo Pedroso <paoloapedroso@gmail.com>
     *
     * @license Apache 2.0
     *
    */

module instr_mem #() ();

endmodule
